library verilog;
use verilog.vl_types.all;
entity tb_lab1 is
end tb_lab1;
